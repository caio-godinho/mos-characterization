** sch_path: /home/caio-godinho/repos/mos-characteriazation/pmos/test_bench.sch
**.subckt test_bench VD VS VB
*.ipin VD
*.ipin VS
*.ipin VB
XM2 net1 net1 VS VB sky130_fd_pr__pfet_g5v0d10v5 L=54.1 W=0.42 nf=1 ad='int((1 + 1)/2) * 0.42 / 1 * 0.29' as='int((1 + 2)/2) * 0.42 / 1 * 0.29'
+ pd='2*int((1 + 1)/2) * (0.42 / 1 + 0.29)' ps='2*int((1 + 2)/2) * (0.42 / 1 + 0.29)' nrd='0.29 / 0.42 ' nrs='0.29 / 0.42 ' sa=0 sb=0
+ sd=0 mult=1 m=1
XM1 VD VD net1 VB sky130_fd_pr__pfet_g5v0d10v5 L=54.1 W=0.42 nf=1 ad='int((1 + 1)/2) * 0.42 / 1 * 0.29' as='int((1 + 2)/2) * 0.42 / 1 * 0.29'
+ pd='2*int((1 + 1)/2) * (0.42 / 1 + 0.29)' ps='2*int((1 + 2)/2) * (0.42 / 1 + 0.29)' nrd='0.29 / 0.42 ' nrs='0.29 / 0.42 ' sa=0 sb=0
+ sd=0 mult=1 m=1
**.ends
.end
