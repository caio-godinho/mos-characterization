********* SIM **********
.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include nmos_characterization.spice

*Vds VD VS 1.5V
Vdgnd VD GND 300mV
*Vgs VG VS 850mV
Vggnd VG GND 850mV
*Vgd VG VD 0.0V
*Vsb VS VB 0.0V
Vbgnd VB GND 0.0V
Vsgnd VS GND 0.0V

.op
*.dc Vgs 0.0 1.5 0.001
*.dc Vds 0.0 3.3 0.01
*.dc Vsb 0.0 1.95 0.01

.control
    setplot new
    setplot const
    let start_l = 0.4
    let stop_l = 0.35
    let delta_l = 0.01
    let l_act = start_l
    let count = 0
    set output_plot = 'unknown1'
    * loop
    while const.l_act le const.stop_l
	let count = $&count + 1
	*alter @m.xm1.msky130_fd_pr__nfet_g5v0d10v5[l] const.l_act
	alter @m.xm1.msky130_fd_pr__nfet_01v8[l] const.l_act
	*save all @m.xm1.msky130_fd_pr__nfet_g5v0d10v5[l] @m.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth]
	save all @m.xm1.msky130_fd_pr__nfet_01v8[l] @m.xm1.msky130_fd_pr__nfet_01v8[vth]
    	run
	*let ids = -I(Vds)
	setplot $output_plot
	*let ids_{$&const.l_act} = dc{$&count}.ids
    	let const.l_act = const.l_act + const.delta_l
	*print @m.xm1.msky130_fd_pr__nfet_g5v0d10v5[vth]
    end
    
    setplot $output_plot
    *plot all vs $&"dc1.v-sweep" ylabel 'Ids' xlabel 'Vds'
    *plot all vs $&"dc1.v-sweep" ylabel 'Ids' xlabel 'Vgs'
    print all.vdgnd#branch all.@m.xm1.msky130_fd_pr__nfet_01v8[vth]
.endc

.end
